---------------------------------------------------------------------------------
library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE WORK.EthConstants.ALL;
---------------------------------------------------------------------------------
ENTITY TxDataState IS
   PORT(
      COUNT_IN : in INTEGER := 0;
      TXD : OUT STD_LOGIC_VECTOR(3 downto 0) := "ZZZZ"
      );
END TxDataState;

---------------------------------------------------------------------------------

ARCHITECTURE Behavioral OF TxDataState IS
BEGIN
   WITH COUNT_IN SELECT
      TXD <= MAC_DESTADDR1 WHEN ETH_DESTADDR1,
             MAC_DESTADDR2 WHEN ETH_DESTADDR2,
             MAC_DESTADDR3 WHEN ETH_DESTADDR3,
             MAC_DESTADDR4 WHEN ETH_DESTADDR4,
             MAC_DESTADDR5 WHEN ETH_DESTADDR5,
             MAC_DESTADDR6 WHEN ETH_DESTADDR6,
             MAC_DESTADDR7 WHEN ETH_DESTADDR7,
             MAC_DESTADDR8 WHEN ETH_DESTADDR8,
             MAC_DESTADDR9 WHEN ETH_DESTADDR9,
             MAC_DESTADDR10 WHEN ETH_DESTADDR10,
             MAC_DESTADDR11 WHEN ETH_DESTADDR11,
             MAC_DESTADDR12 WHEN ETH_DESTADDR12,
             MAC_SRCADDR1 WHEN ETH_SRCADDR1,
             MAC_SRCADDR2 WHEN ETH_SRCADDR2,
             MAC_SRCADDR3 WHEN ETH_SRCADDR3,
             MAC_SRCADDR4 WHEN ETH_SRCADDR4,
             MAC_SRCADDR5 WHEN ETH_SRCADDR5,
             MAC_SRCADDR6 WHEN ETH_SRCADDR6,
             MAC_SRCADDR7 WHEN ETH_SRCADDR7,
             MAC_SRCADDR8 WHEN ETH_SRCADDR8,
             MAC_SRCADDR9 WHEN ETH_SRCADDR9,
             MAC_SRCADDR10 WHEN ETH_SRCADDR10,
             MAC_SRCADDR11 WHEN ETH_SRCADDR11,
             MAC_SRCADDR12 WHEN ETH_SRCADDR12,
             ETHERTYPE1 WHEN ETH_TYPE1,
             ETHERTYPE2 WHEN ETH_TYPE2,
             ETHERTYPE3 WHEN ETH_TYPE3,
             ETHERTYPE4 WHEN ETH_TYPE4,
             IP_VER WHEN ETH_IPV4_IHL,
             IP_IHL WHEN ETH_IPV4_VER,
             IP_SRVTP1 WHEN ETH_IPV4_SRVTP1,
             IP_SRVTP2 WHEN ETH_IPV4_SRVTP2,
             IP_LENG1 WHEN ETH_IPV4_LNG1,
             IP_LENG2 WHEN ETH_IPV4_LNG2,
             IP_LENG3 WHEN ETH_IPV4_LNG3,
             IP_LENG4 WHEN ETH_IPV4_LNG4,
             IP_ID WHEN ETH_IPV4_ID1,
             IP_ID WHEN ETH_IPV4_ID2,
             IP_ID WHEN ETH_IPV4_ID3,
             IP_ID WHEN ETH_IPV4_ID4,
             IP_FLAGS WHEN ETH_IPV4_FLG,
             IP_OFFSET0 WHEN ETH_IPV4_FRAGOFF1,
             IP_OFFSET1 WHEN ETH_IPV4_FRAGOFF2,
             IP_OFFSET2 WHEN ETH_IPV4_FRAGOFF3,
             IP_TTL1 WHEN ETH_IPV4_LIVETIME1,
             IP_TTL2 WHEN ETH_IPV4_LIVETIME2,
             IP_PROTOCOL1 WHEN ETH_IPV4_PROTOCOL1,
             IP_PROTOCOL2 WHEN ETH_IPV4_PROTOCOL2,
             IP_HDCHKSUM1 WHEN ETH_IPV4_HEADERCHKSM1,
             IP_HDCHKSUM2 WHEN ETH_IPV4_HEADERCHKSM2,
             IP_HDCHKSUM3 WHEN ETH_IPV4_HEADERCHKSM3,
             IP_HDCHKSUM4 WHEN ETH_IPV4_HEADERCHKSM4,
             IP_SRCIP1 WHEN ETH_IPV4_SRCIP1,
             IP_SRCIP2 WHEN ETH_IPV4_SRCIP2,
             IP_SRCIP3 WHEN ETH_IPV4_SRCIP3,
             IP_SRCIP4 WHEN ETH_IPV4_SRCIP4,
             IP_SRCIP5 WHEN ETH_IPV4_SRCIP5,
             IP_SRCIP6 WHEN ETH_IPV4_SRCIP6,
             IP_SRCIP7 WHEN ETH_IPV4_SRCIP7,
             IP_SRCIP8 WHEN ETH_IPV4_SRCIP8,
             IP_DSTIP1 WHEN ETH_IPV4_DSTIP1,
             IP_DSTIP2 WHEN ETH_IPV4_DSTIP2,
             IP_DSTIP3 WHEN ETH_IPV4_DSTIP3,
             IP_DSTIP4 WHEN ETH_IPV4_DSTIP4,
             IP_DSTIP5 WHEN ETH_IPV4_DSTIP5,
             IP_DSTIP6 WHEN ETH_IPV4_DSTIP6,
             IP_DSTIP7 WHEN ETH_IPV4_DSTIP7,
             IP_DSTIP8 WHEN ETH_IPV4_DSTIP8,
             UDP_SRCADR1 WHEN ETH_IPV4_UDP_SRCADR1,
             UDP_SRCADR2 WHEN ETH_IPV4_UDP_SRCADR2,
             UDP_SRCADR3 WHEN ETH_IPV4_UDP_SRCADR3,
             UDP_SRCADR4 WHEN ETH_IPV4_UDP_SRCADR4,
             UDP_DSTADR1 WHEN ETH_IPV4_UDP_DSTADR1,
             UDP_DSTADR2 WHEN ETH_IPV4_UDP_DSTADR2,
             UDP_DSTADR3 WHEN ETH_IPV4_UDP_DSTADR3,
             UDP_DSTADR4 WHEN ETH_IPV4_UDP_DSTADR4,
             UDP_LENG1 WHEN ETH_IPV4_UDP_LENG1,
             UDP_LENG2 WHEN ETH_IPV4_UDP_LENG2,
             UDP_LENG3 WHEN ETH_IPV4_UDP_LENG3,
             UDP_LENG4 WHEN ETH_IPV4_UDP_LENG4,
             UDP_CHKSUM0 WHEN ETH_IPV4_UDP_CHKSUM1,
             UDP_CHKSUM1 WHEN ETH_IPV4_UDP_CHKSUM2,
             UDP_CHKSUM2 WHEN ETH_IPV4_UDP_CHKSUM3,
             UDP_CHKSUM3 WHEN ETH_IPV4_UDP_CHKSUM4,
             
             --
             -- Need to input camera data here
             --
             
             "ZZZZ" WHEN OTHERS;

---------------------------------------------------------------------------------
END Behavioral;
