--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

package EthConstants is

-- type <new_type> is
--  record
--    <type_name>        : std_logic_vector( 7 downto 0);
--    <type_name>        : std_logic;
-- end record;
--
-- Declare constants
--
CONSTANT ETH_SFD1 : INTEGER := 11;
CONSTANT ETH_SFD2 : INTEGER := ETH_SFD1 + 1;
CONSTANT ETH_DESTADDR2 : INTEGER := ETH_SFD2 + 1;
CONSTANT ETH_DESTADDR1 : INTEGER := ETH_DESTADDR2 + 1;
CONSTANT ETH_DESTADDR4 : INTEGER := ETH_DESTADDR1 + 1;
CONSTANT ETH_DESTADDR3 : INTEGER := ETH_DESTADDR4 + 1;
CONSTANT ETH_DESTADDR6 : INTEGER := ETH_DESTADDR3 + 1;
CONSTANT ETH_DESTADDR5 : INTEGER := ETH_DESTADDR6 + 1;
CONSTANT ETH_DESTADDR8 : INTEGER := ETH_DESTADDR5 + 1;
CONSTANT ETH_DESTADDR7 : INTEGER := ETH_DESTADDR8 + 1;
CONSTANT ETH_DESTADDR10 : INTEGER := ETH_DESTADDR7 + 1;
CONSTANT ETH_DESTADDR9 : INTEGER := ETH_DESTADDR10 + 1;
CONSTANT ETH_DESTADDR12 : INTEGER := ETH_DESTADDR9 + 1;
CONSTANT ETH_DESTADDR11 : INTEGER := ETH_DESTADDR12 + 1;
CONSTANT ETH_SRCADDR2 : INTEGER := ETH_DESTADDR11 + 1;
CONSTANT ETH_SRCADDR1 : INTEGER := ETH_SRCADDR2 + 1;
CONSTANT ETH_SRCADDR4 : INTEGER := ETH_SRCADDR1 + 1;
CONSTANT ETH_SRCADDR3 : INTEGER := ETH_SRCADDR4 + 1;
CONSTANT ETH_SRCADDR6 : INTEGER := ETH_SRCADDR3 + 1;
CONSTANT ETH_SRCADDR5 : INTEGER := ETH_SRCADDR6 + 1;
CONSTANT ETH_SRCADDR8 : INTEGER := ETH_SRCADDR5 + 1;
CONSTANT ETH_SRCADDR7 : INTEGER := ETH_SRCADDR8 + 1;
CONSTANT ETH_SRCADDR10 : INTEGER := ETH_SRCADDR7 + 1;
CONSTANT ETH_SRCADDR9 : INTEGER := ETH_SRCADDR10 + 1;
CONSTANT ETH_SRCADDR12 : INTEGER := ETH_SRCADDR9 + 1;
CONSTANT ETH_SRCADDR11 : INTEGER := ETH_SRCADDR12 + 1;
CONSTANT ETH_TYPE2 : INTEGER := ETH_SRCADDR11 + 1;
CONSTANT ETH_TYPE1 : INTEGER := ETH_TYPE2 + 1;
CONSTANT ETH_TYPE4 : INTEGER := ETH_TYPE1 + 1;
CONSTANT ETH_TYPE3 : INTEGER := ETH_TYPE4 + 1;


-- IPv4 Header Offsets

-- 20Bytes
-- 0  |0____.____|1____.____|2____.____|3____.____|
-- 4  | Ver |Leng|Serv Type |     Total Length    |
-- 8  |    Identification   |Flags|Fragment Offset|
-- 12 |    TTL   | Protocol | Header Checksum     |
-- 16 |             Source Address                |
-- 20 |            Destination Address            |

CONSTANT ETH_IPV4_IHL : INTEGER := ETH_TYPE3 + 1;
CONSTANT ETH_IPV4_VER : INTEGER := ETH_IPV4_IHL + 1;
CONSTANT ETH_IPV4_SRVTP2 : INTEGER := ETH_IPV4_VER + 1;
CONSTANT ETH_IPV4_SRVTP1 : INTEGER := ETH_IPV4_SRVTP2 + 1;
CONSTANT ETH_IPV4_LNG2 : INTEGER := ETH_IPV4_SRVTP1 + 1;
CONSTANT ETH_IPV4_LNG1 : INTEGER := ETH_IPV4_LNG2 + 1;
CONSTANT ETH_IPV4_LNG4 : INTEGER := ETH_IPV4_LNG1 + 1;
CONSTANT ETH_IPV4_LNG3 : INTEGER := ETH_IPV4_LNG4 + 1;
CONSTANT ETH_IPV4_ID2 : INTEGER := ETH_IPV4_LNG3 + 1;
CONSTANT ETH_IPV4_ID1 : INTEGER := ETH_IPV4_ID2 + 1;
CONSTANT ETH_IPV4_ID4 : INTEGER := ETH_IPV4_ID1 + 1;
CONSTANT ETH_IPV4_ID3 : INTEGER := ETH_IPV4_ID4 + 1;
CONSTANT ETH_IPV4_FRAGOFF1 : INTEGER := ETH_IPV4_ID3 + 1;
CONSTANT ETH_IPV4_FLG : INTEGER := ETH_IPV4_FRAGOFF1 + 1;
CONSTANT ETH_IPV4_FRAGOFF3 : INTEGER := ETH_IPV4_FLG + 1;
CONSTANT ETH_IPV4_FRAGOFF2 : INTEGER := ETH_IPV4_FRAGOFF3 + 1;
CONSTANT ETH_IPV4_LIVETIME2 : INTEGER := ETH_IPV4_FRAGOFF2 + 1;
CONSTANT ETH_IPV4_LIVETIME1 : INTEGER := ETH_IPV4_LIVETIME2 + 1;
CONSTANT ETH_IPV4_PROTOCOL2 : INTEGER := ETH_IPV4_LIVETIME1 + 1;
CONSTANT ETH_IPV4_PROTOCOL1 : INTEGER := ETH_IPV4_PROTOCOL2 + 1;
CONSTANT ETH_IPV4_HEADERCHKSM2 : INTEGER := ETH_IPV4_PROTOCOL1 + 1;
CONSTANT ETH_IPV4_HEADERCHKSM1 : INTEGER := ETH_IPV4_HEADERCHKSM2 + 1;
CONSTANT ETH_IPV4_HEADERCHKSM4 : INTEGER := ETH_IPV4_HEADERCHKSM1 + 1;
CONSTANT ETH_IPV4_HEADERCHKSM3 : INTEGER := ETH_IPV4_HEADERCHKSM4 + 1;
CONSTANT ETH_IPV4_SRCIP2 : INTEGER := ETH_IPV4_HEADERCHKSM3 + 1;
CONSTANT ETH_IPV4_SRCIP1 : INTEGER := ETH_IPV4_SRCIP2 + 1;
CONSTANT ETH_IPV4_SRCIP4 : INTEGER := ETH_IPV4_SRCIP1 + 1;
CONSTANT ETH_IPV4_SRCIP3 : INTEGER := ETH_IPV4_SRCIP4 + 1;
CONSTANT ETH_IPV4_SRCIP6 : INTEGER := ETH_IPV4_SRCIP3 + 1;
CONSTANT ETH_IPV4_SRCIP5 : INTEGER := ETH_IPV4_SRCIP6 + 1;
CONSTANT ETH_IPV4_SRCIP8 : INTEGER := ETH_IPV4_SRCIP5 + 1;
CONSTANT ETH_IPV4_SRCIP7 : INTEGER := ETH_IPV4_SRCIP8 + 1;
CONSTANT ETH_IPV4_DSTIP2 : INTEGER := ETH_IPV4_SRCIP7 + 1;
CONSTANT ETH_IPV4_DSTIP1 : INTEGER := ETH_IPV4_DSTIP2 + 1;
CONSTANT ETH_IPV4_DSTIP4 : INTEGER := ETH_IPV4_DSTIP1 + 1;
CONSTANT ETH_IPV4_DSTIP3 : INTEGER := ETH_IPV4_DSTIP4 + 1;
CONSTANT ETH_IPV4_DSTIP6 : INTEGER := ETH_IPV4_DSTIP3 + 1;
CONSTANT ETH_IPV4_DSTIP5 : INTEGER := ETH_IPV4_DSTIP6 + 1;
CONSTANT ETH_IPV4_DSTIP8 : INTEGER := ETH_IPV4_DSTIP5 + 1;
CONSTANT ETH_IPV4_DSTIP7 : INTEGER := ETH_IPV4_DSTIP8 + 1;
CONSTANT ETH_IPV4_PAYLOAD : INTEGER := ETH_IPV4_DSTIP7 + 1;


-- UDP Header Offsets
-- 8Bytes
-- 0  |0____.____|1____.____|2____.____|3____.____|
-- 4  |    Source Address   | Destination Address |
-- 8  |        Length       |       Checksum      |
CONSTANT ETH_IPV4_UDP_SRCADR2 : INTEGER := ETH_IPV4_DSTIP7 + 1;
CONSTANT ETH_IPV4_UDP_SRCADR1 : INTEGER := ETH_IPV4_UDP_SRCADR2 + 1;
CONSTANT ETH_IPV4_UDP_SRCADR4 : INTEGER := ETH_IPV4_UDP_SRCADR1 + 1;
CONSTANT ETH_IPV4_UDP_SRCADR3 : INTEGER := ETH_IPV4_UDP_SRCADR4 + 1;
CONSTANT ETH_IPV4_UDP_DSTADR2 : INTEGER := ETH_IPV4_UDP_SRCADR3 + 1;
CONSTANT ETH_IPV4_UDP_DSTADR1 : INTEGER := ETH_IPV4_UDP_DSTADR2 + 1;
CONSTANT ETH_IPV4_UDP_DSTADR4 : INTEGER := ETH_IPV4_UDP_DSTADR1 + 1;
CONSTANT ETH_IPV4_UDP_DSTADR3 : INTEGER := ETH_IPV4_UDP_DSTADR4 + 1;
CONSTANT ETH_IPV4_UDP_LENG2 : INTEGER   := ETH_IPV4_UDP_DSTADR3 + 1;
CONSTANT ETH_IPV4_UDP_LENG1 : INTEGER   := ETH_IPV4_UDP_LENG2 + 1;
CONSTANT ETH_IPV4_UDP_LENG4 : INTEGER   := ETH_IPV4_UDP_LENG1 + 1;
CONSTANT ETH_IPV4_UDP_LENG3 : INTEGER   := ETH_IPV4_UDP_LENG4 + 1;
CONSTANT ETH_IPV4_UDP_CHKSUM2 : INTEGER := ETH_IPV4_UDP_LENG3 + 1;
CONSTANT ETH_IPV4_UDP_CHKSUM1 : INTEGER := ETH_IPV4_UDP_CHKSUM2 + 1;
CONSTANT ETH_IPV4_UDP_CHKSUM4 : INTEGER := ETH_IPV4_UDP_CHKSUM1 + 1;
CONSTANT ETH_IPV4_UDP_CHKSUM3 : INTEGER := ETH_IPV4_UDP_CHKSUM4 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N2 : INTEGER := ETH_IPV4_UDP_CHKSUM3 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N1 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N2 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N4 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N1  + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N3 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N4 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N6 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N3 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N5 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N6 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N8 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N5 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N7 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N8 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N10 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N7 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N9 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N10 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N12 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N9 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N11 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N12 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N14 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N11 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N13 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N14 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N16 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N13 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N15 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N16 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N18 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N15 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N17 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N18 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N20 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N17 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N19 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N20 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N22 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N19 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N21 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N22 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N24 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N21 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N23 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N24 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N26 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N23 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N25 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N26 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N28 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N25 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N27 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N28 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N30 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N27 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N29 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N30 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N32 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N29 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N31 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N32 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N34 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N31 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N33 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N34 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N36 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N33 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N35 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N36 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N38 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N35 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N37 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N38 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N40 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N37 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N39 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N40 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N42 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N39 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N41 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N42 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N44 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N41 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N43 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N44 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N46 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N43 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N45 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N46 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N48 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N45 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD_N47 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N48 + 1;
CONSTANT ETH_IPV4_UDP_PAYLOAD : INTEGER := ETH_IPV4_UDP_PAYLOAD_N47;


CONSTANT ETH_IPV4_UDP_ENDOFPAYLOAD : INTEGER := ETH_IPV4_UDP_PAYLOAD; -- = (ETH_IPV4_UDP_PAYLOAD) + (UDP Payload size)
CONSTANT ETH_IP_ENDOFPAYLOAD : INTEGER := ETH_IPV4_UDP_PAYLOAD; -- = (ETH_IPV4_UDP_PAYLOAD) + (UDP Payload size)
CONSTANT ETH_PAYLOAD : INTEGER := ETH_IPV4_UDP_PAYLOAD; -- Consider changing this to where CRC begins

CONSTANT ETH_CRC2 : INTEGER := ETH_IPV4_UDP_PAYLOAD + 1;
CONSTANT ETH_CRC1 : INTEGER := ETH_CRC2 + 1;
CONSTANT ETH_CRC4 : INTEGER := ETH_CRC1 + 1;
CONSTANT ETH_CRC3 : INTEGER := ETH_CRC4 + 1;
CONSTANT ETH_CRC6 : INTEGER := ETH_CRC3 + 1;
CONSTANT ETH_CRC5 : INTEGER := ETH_CRC6 + 1;
CONSTANT ETH_CRC8 : INTEGER := ETH_CRC5 + 1;
CONSTANT ETH_CRC7 : INTEGER := ETH_CRC8 + 1;

CONSTANT ETH_END_FRAME : INTEGER := ETH_CRC7 + 1;



CONSTANT CRC_ETHERNETCOUNT3 : INTEGER := 1;
CONSTANT CRC_ETHERNETCOUNT4 : INTEGER := CRC_ETHERNETCOUNT3 + 1;
CONSTANT CRC_ETHERNETCOUNT5 : INTEGER := CRC_ETHERNETCOUNT4 + 1;
CONSTANT CRC_ETHERNETCOUNT6 : INTEGER := CRC_ETHERNETCOUNT5 + 1;
CONSTANT CRC_ETHERNETCOUNT7 : INTEGER := CRC_ETHERNETCOUNT6 + 1;
CONSTANT CRC_ETHERNETCOUNT8 : INTEGER := CRC_ETHERNETCOUNT7 + 1;
CONSTANT CRC_ETHERNETCOUNT9 : INTEGER := CRC_ETHERNETCOUNT8 + 1;
CONSTANT CRC_ETHERNETCOUNT10 : INTEGER := CRC_ETHERNETCOUNT9 + 1;
CONSTANT CRC_ETHERNETCOUNT11 : INTEGER := CRC_ETHERNETCOUNT10 + 1;
CONSTANT CRC_ETHERNETCOUNT12 : INTEGER := CRC_ETHERNETCOUNT11 + 1;
CONSTANT CRC_ETHERNETCOUNT13 : INTEGER := CRC_ETHERNETCOUNT12 + 1;
CONSTANT CRC_ETHERNETCOUNT14 : INTEGER := CRC_ETHERNETCOUNT13 + 1;
CONSTANT CRC_ETHERNETCOUNT15 : INTEGER := CRC_ETHERNETCOUNT14 + 1;
CONSTANT CRC_ETHERNETCOUNT16 : INTEGER := CRC_ETHERNETCOUNT15 + 1;
CONSTANT CRC_ETHERNETCOUNT17 : INTEGER := CRC_ETHERNETCOUNT16 + 1;
CONSTANT CRC_ETHERNETCOUNT18 : INTEGER := CRC_ETHERNETCOUNT17 + 1;
CONSTANT CRC_ETHERNETCOUNT19 : INTEGER := CRC_ETHERNETCOUNT18 + 1;
CONSTANT CRC_ETHERNETCOUNT20 : INTEGER := CRC_ETHERNETCOUNT19 + 1;
CONSTANT CRC_ETHERNETCOUNT21 : INTEGER := CRC_ETHERNETCOUNT20 + 1;
CONSTANT CRC_ETHERNETCOUNT22 : INTEGER := CRC_ETHERNETCOUNT21 + 1;
CONSTANT CRC_ETHERNETCOUNT23 : INTEGER := CRC_ETHERNETCOUNT22 + 1;
CONSTANT CRC_ETHERNETCOUNT24 : INTEGER := CRC_ETHERNETCOUNT23 + 1;
CONSTANT CRC_ETHERNETCOUNT25 : INTEGER := CRC_ETHERNETCOUNT24 + 1;
CONSTANT CRC_ETHERNETCOUNT26 : INTEGER := CRC_ETHERNETCOUNT25 + 1;
CONSTANT CRC_ETHERNETCOUNT27 : INTEGER := CRC_ETHERNETCOUNT26 + 1;
CONSTANT CRC_ETHERNETCOUNT28 : INTEGER := CRC_ETHERNETCOUNT27 + 1;
CONSTANT CRC_ETHERNETCOUNT29 : INTEGER := CRC_ETHERNETCOUNT28 + 1;
CONSTANT CRC_ETHERNETCOUNT30 : INTEGER := CRC_ETHERNETCOUNT29 + 1;
CONSTANT CRC_ETHERNETCOUNT31 : INTEGER := CRC_ETHERNETCOUNT30 + 1;
CONSTANT CRC_ETHERNETCOUNT32 : INTEGER := CRC_ETHERNETCOUNT31 + 1;
CONSTANT CRC_ETHERNETCOUNT33 : INTEGER := CRC_ETHERNETCOUNT32 + 1;
CONSTANT CRC_ETHERNETCOUNT34 : INTEGER := CRC_ETHERNETCOUNT33 + 1;
CONSTANT CRC_ETHERNETCOUNT35 : INTEGER := CRC_ETHERNETCOUNT34 + 1;
CONSTANT CRC_ETHERNETCOUNT36 : INTEGER := CRC_ETHERNETCOUNT35 + 1;
CONSTANT CRC_ETHERNETCOUNT37 : INTEGER := CRC_ETHERNETCOUNT36 + 1;
CONSTANT CRC_ETHERNETCOUNT38 : INTEGER := CRC_ETHERNETCOUNT37 + 1;
CONSTANT CRC_ETHERNETCOUNT39 : INTEGER := CRC_ETHERNETCOUNT38 + 1;
CONSTANT CRC_ETHERNETCOUNT40 : INTEGER := CRC_ETHERNETCOUNT39 + 1;
CONSTANT CRC_ETHERNETCOUNT41 : INTEGER := CRC_ETHERNETCOUNT40 + 1;
CONSTANT CRC_ETHERNETCOUNT42 : INTEGER := CRC_ETHERNETCOUNT41 + 1;
CONSTANT CRC_ETHERNETCOUNT43 : INTEGER := CRC_ETHERNETCOUNT42 + 1;
CONSTANT CRC_ETHERNETCOUNT44 : INTEGER := CRC_ETHERNETCOUNT43 + 1;
CONSTANT CRC_ETHERNETCOUNT45 : INTEGER := CRC_ETHERNETCOUNT44 + 1;
CONSTANT CRC_ETHERNETCOUNT46 : INTEGER := CRC_ETHERNETCOUNT45 + 1;
CONSTANT CRC_ETHERNETCOUNT47 : INTEGER := CRC_ETHERNETCOUNT46 + 1;
CONSTANT CRC_ETHERNETCOUNT48 : INTEGER := CRC_ETHERNETCOUNT47 + 1;
CONSTANT CRC_ETHERNETCOUNT49 : INTEGER := CRC_ETHERNETCOUNT48 + 1;
CONSTANT CRC_ETHERNETCOUNT50 : INTEGER := CRC_ETHERNETCOUNT49 + 1;
CONSTANT CRC_ETHERNETCOUNT51 : INTEGER := CRC_ETHERNETCOUNT50 + 1;
CONSTANT CRC_ETHERNETCOUNT52 : INTEGER := CRC_ETHERNETCOUNT51 + 1;
CONSTANT CRC_ETHERNETCOUNT53 : INTEGER := CRC_ETHERNETCOUNT52 + 1;
CONSTANT CRC_ETHERNETCOUNT54 : INTEGER := CRC_ETHERNETCOUNT53 + 1;
CONSTANT CRC_ETHERNETCOUNT55 : INTEGER := CRC_ETHERNETCOUNT54 + 1;
CONSTANT CRC_ETHERNETCOUNT56 : INTEGER := CRC_ETHERNETCOUNT55 + 1;
CONSTANT CRC_ETHERNETCOUNT57 : INTEGER := CRC_ETHERNETCOUNT56 + 1;
CONSTANT CRC_ETHERNETCOUNT58 : INTEGER := CRC_ETHERNETCOUNT57 + 1;
CONSTANT CRC_ETHERNETCOUNT59 : INTEGER := CRC_ETHERNETCOUNT58 + 1;
CONSTANT CRC_ETHERNETCOUNT60 : INTEGER := CRC_ETHERNETCOUNT59 + 1;
CONSTANT CRC_ETHERNETCOUNT61 : INTEGER := CRC_ETHERNETCOUNT60 + 1;
CONSTANT CRC_ETHERNETCOUNT62 : INTEGER := CRC_ETHERNETCOUNT61 + 1;
CONSTANT CRC_ETHERNETCOUNT63 : INTEGER := CRC_ETHERNETCOUNT62 + 1;
CONSTANT CRC_ETHERNETCOUNT64 : INTEGER := CRC_ETHERNETCOUNT63 + 1;
CONSTANT CRC_ETHERNETCOUNT65 : INTEGER := CRC_ETHERNETCOUNT64 + 1;
CONSTANT CRC_ETHERNETCOUNT66 : INTEGER := CRC_ETHERNETCOUNT65 + 1;
CONSTANT CRC_ETHERNETCOUNT67 : INTEGER := CRC_ETHERNETCOUNT66 + 1;
CONSTANT CRC_ETHERNETCOUNT68 : INTEGER := CRC_ETHERNETCOUNT67 + 1;
CONSTANT CRC_ETHERNETCOUNT69 : INTEGER := CRC_ETHERNETCOUNT68 + 1;











--------------------------------------------------------------------------------
-- Defined Values

CONSTANT ETH_FRAMEGAP : INTEGER := ETH_CRC7 + 24;
CONSTANT ETHPREAMBLE : STD_LOGIC_VECTOR := "1010";
CONSTANT SFD1 : STD_LOGIC_VECTOR(7 downto 0) := X"05";
CONSTANT SFD2 : STD_LOGIC_VECTOR(7 downto 0) := X"0D";
CONSTANT BROADCAST : STD_LOGIC_VECTOR(7 downto 0) := X"0F";
CONSTANT MAC_DESTADDR1 : STD_LOGIC_VECTOR(7 downto 0) := X"00";  -- 0 -- 00-1d-92-f3-31-53
CONSTANT MAC_DESTADDR2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";  -- 0
CONSTANT MAC_DESTADDR3 : STD_LOGIC_VECTOR(7 downto 0) := X"01";  -- 1
CONSTANT MAC_DESTADDR4 : STD_LOGIC_VECTOR(7 downto 0) := X"0D";  -- D
CONSTANT MAC_DESTADDR5 : STD_LOGIC_VECTOR(7 downto 0) := X"09";  -- 9
CONSTANT MAC_DESTADDR6 : STD_LOGIC_VECTOR(7 downto 0) := X"02";  -- 2
CONSTANT MAC_DESTADDR7 : STD_LOGIC_VECTOR(7 downto 0) := X"0F";  -- F
CONSTANT MAC_DESTADDR8 : STD_LOGIC_VECTOR(7 downto 0) := X"03";  -- 3
CONSTANT MAC_DESTADDR9 : STD_LOGIC_VECTOR(7 downto 0) := X"03";  -- 3
CONSTANT MAC_DESTADDR10 : STD_LOGIC_VECTOR(7 downto 0) := X"01";  -- 1
CONSTANT MAC_DESTADDR11 : STD_LOGIC_VECTOR(7 downto 0) := X"05";  -- 5
CONSTANT MAC_DESTADDR12 : STD_LOGIC_VECTOR(7 downto 0) := X"03";  -- 3
CONSTANT MAC_SRCADDR1 : STD_LOGIC_VECTOR(7 downto 0) := X"0A";  -- A -- A3-1C-6D-DF-B6-B6
CONSTANT MAC_SRCADDR2 : STD_LOGIC_VECTOR(7 downto 0) := X"03";  -- 3
CONSTANT MAC_SRCADDR3 : STD_LOGIC_VECTOR(7 downto 0) := X"01";  -- 1
CONSTANT MAC_SRCADDR4 : STD_LOGIC_VECTOR(7 downto 0) := X"0C";  -- C
CONSTANT MAC_SRCADDR5 : STD_LOGIC_VECTOR(7 downto 0) := X"06";  -- 6
CONSTANT MAC_SRCADDR6 : STD_LOGIC_VECTOR(7 downto 0) := X"0D";  -- D
CONSTANT MAC_SRCADDR7 : STD_LOGIC_VECTOR(7 downto 0) := X"0D";  -- D
CONSTANT MAC_SRCADDR8 : STD_LOGIC_VECTOR(7 downto 0) := X"0F";  -- F
CONSTANT MAC_SRCADDR9 : STD_LOGIC_VECTOR(7 downto 0) := X"0B";  -- B
CONSTANT MAC_SRCADDR10 : STD_LOGIC_VECTOR(7 downto 0) := X"06"; -- 6
CONSTANT MAC_SRCADDR11 : STD_LOGIC_VECTOR(7 downto 0) := X"0B"; -- B
CONSTANT MAC_SRCADDR12 : STD_LOGIC_VECTOR(7 downto 0) := X"06"; -- 6
CONSTANT ETHERTYPE1 : STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- 0
CONSTANT ETHERTYPE2 : STD_LOGIC_VECTOR(7 downto 0) := X"08"; -- 8
CONSTANT ETHERTYPE3 : STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- 0
CONSTANT ETHERTYPE4 : STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- 0
CONSTANT CRC1 : STD_LOGIC_VECTOR(7 downto 0) := X"07"; -- bd890fc8 --> http://www.zorc.breitbandkatze.de/crc.html
CONSTANT CRC2 : STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- d6fe9a4b --> Test bench
CONSTANT CRC3 : STD_LOGIC_VECTOR(7 downto 0) := X"07";
CONSTANT CRC4 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT CRC5 : STD_LOGIC_VECTOR(7 downto 0) := X"0A";
CONSTANT CRC6 : STD_LOGIC_VECTOR(7 downto 0) := X"0D";
CONSTANT CRC7 : STD_LOGIC_VECTOR(7 downto 0) := X"0F";
CONSTANT CRC8 : STD_LOGIC_VECTOR(7 downto 0) := X"0C";

-- IPv4 Header Constants
CONSTANT IP_VER : STD_LOGIC_VECTOR(7 downto 0) := X"04";
CONSTANT IP_IHL : STD_LOGIC_VECTOR(7 downto 0) := X"05";
CONSTANT IP_SRVTP1 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_SRVTP2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_LENG1 : STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- = (20 Byte IP header) + (8 Byte UDP header) + (24 Byte UDP payload) = 52
CONSTANT IP_LENG2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_LENG3 : STD_LOGIC_VECTOR(7 downto 0) := X"03";
CONSTANT IP_LENG4 : STD_LOGIC_VECTOR(7 downto 0) := X"04";
CONSTANT IP_ID0 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_ID1 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_FLAGS : STD_LOGIC_VECTOR(7 downto 0) := X"04"; -- 11:7
CONSTANT IP_OFFSET0: STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_OFFSET1: STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_OFFSET2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_TTL1 : STD_LOGIC_VECTOR(7 downto 0) := X"0F";
CONSTANT IP_TTL2 : STD_LOGIC_VECTOR(7 downto 0) := X"0F";
CONSTANT IP_PROTOCOL1 : STD_LOGIC_VECTOR(7 downto 0) := X"01"; -- UDP Protocol ID
CONSTANT IP_PROTOCOL2 : STD_LOGIC_VECTOR(7 downto 0) := X"01";
CONSTANT IP_HDCHKSUM1 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_HDCHKSUM2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_HDCHKSUM3 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_HDCHKSUM4 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_SRCIP1 : STD_LOGIC_VECTOR(7 downto 0) := X"0C"; -- IP source is 192
CONSTANT IP_SRCIP2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_SRCIP3 : STD_LOGIC_VECTOR(7 downto 0) := X"0A"; -- .168
CONSTANT IP_SRCIP4 : STD_LOGIC_VECTOR(7 downto 0) := X"08";
CONSTANT IP_SRCIP5 : STD_LOGIC_VECTOR(7 downto 0) := X"08"; -- .137
CONSTANT IP_SRCIP6 : STD_LOGIC_VECTOR(7 downto 0) := X"09";
CONSTANT IP_SRCIP7 : STD_LOGIC_VECTOR(7 downto 0) := X"07"; -- .120
CONSTANT IP_SRCIP8 : STD_LOGIC_VECTOR(7 downto 0) := X"08";
CONSTANT IP_DSTIP1 : STD_LOGIC_VECTOR(7 downto 0) := X"0C"; -- IP destination is 192
CONSTANT IP_DSTIP2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT IP_DSTIP3 : STD_LOGIC_VECTOR(7 downto 0) := X"0A"; -- .168
CONSTANT IP_DSTIP4 : STD_LOGIC_VECTOR(7 downto 0) := X"08";
CONSTANT IP_DSTIP5 : STD_LOGIC_VECTOR(7 downto 0) := X"08"; -- .137
CONSTANT IP_DSTIP6 : STD_LOGIC_VECTOR(7 downto 0) := X"09";
CONSTANT IP_DSTIP7 : STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- .1
CONSTANT IP_DSTIP8 : STD_LOGIC_VECTOR(7 downto 0) := X"01";

-- UDP Header Constants
CONSTANT UDP_SRCADR1 : STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- Least significant nibble
CONSTANT UDP_SRCADR2 : STD_LOGIC_VECTOR(7 downto 0) := X"0A";
CONSTANT UDP_SRCADR3 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT UDP_SRCADR4 : STD_LOGIC_VECTOR(7 downto 0) := X"0A"; -- Most significant nibble
CONSTANT UDP_DSTADR1 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT UDP_DSTADR2 : STD_LOGIC_VECTOR(7 downto 0) := X"0C";
CONSTANT UDP_DSTADR3 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT UDP_DSTADR4 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT UDP_LENG1 : STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- (8Byte header) + (24Byte payload) = 32
CONSTANT UDP_LENG2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT UDP_LENG3 : STD_LOGIC_VECTOR(7 downto 0) := X"02";
CONSTANT UDP_LENG4 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
CONSTANT UDP_CHKSUM0 : STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- 0
CONSTANT UDP_CHKSUM1: STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- 0
CONSTANT UDP_CHKSUM2: STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- 0
CONSTANT UDP_CHKSUM3: STD_LOGIC_VECTOR(7 downto 0) := X"00"; -- 0
CONSTANT UDP_DATA_N1 : STD_LOGIC_VECTOR(7 downto 0) := X"01";
CONSTANT UDP_DATA_N2 : STD_LOGIC_VECTOR(7 downto 0) := X"02";
CONSTANT UDP_DATA_N3 : STD_LOGIC_VECTOR(7 downto 0) := X"03";
CONSTANT UDP_DATA_N4 : STD_LOGIC_VECTOR(7 downto 0) := X"04";
CONSTANT UDP_DATA_N5 : STD_LOGIC_VECTOR(7 downto 0) := X"05";
CONSTANT UDP_DATA_N6 : STD_LOGIC_VECTOR(7 downto 0) := X"06";
CONSTANT UDP_DATA_N7 : STD_LOGIC_VECTOR(7 downto 0) := X"07";
CONSTANT UDP_DATA_N8 : STD_LOGIC_VECTOR(7 downto 0) := X"08";
CONSTANT UDP_DATA_N9 : STD_LOGIC_VECTOR(7 downto 0) := X"09";
CONSTANT UDP_DATA_NA : STD_LOGIC_VECTOR(7 downto 0) := X"0A";
CONSTANT UDP_DATA_NB : STD_LOGIC_VECTOR(7 downto 0) := X"0B";
CONSTANT UDP_DATA_NC : STD_LOGIC_VECTOR(7 downto 0) := X"0C";
CONSTANT UDP_DATA_ND : STD_LOGIC_VECTOR(7 downto 0) := X"0D";
CONSTANT UDP_DATA_NE : STD_LOGIC_VECTOR(7 downto 0) := X"0E";
CONSTANT UDP_DATA_NF : STD_LOGIC_VECTOR(7 downto 0) := X"0F";
CONSTANT UDP_DATA_N0 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
--CONSTANT END_OF_TX1 : STD_LOGIC_VECTOR := "01101";
--CONSTANT END_OF_TX2 : STD_LOGIC_VECTOR := "00111";


---------------------------------------------------------------------------------
-- Declare functions and procedure
--
-- function <function_name>  (signal <signal_name> : in <type_declaration>) return <type_declaration>;
-- procedure <procedure_name> (<type_declaration> <constant_name>	: in <type_declaration>);
--

end EthConstants;

package body EthConstants is

---- Example 1
--  function <function_name>  (signal <signal_name> : in <type_declaration>  ) return <type_declaration> is
--    variable <variable_name>     : <type_declaration>;
--  begin
--    <variable_name> := <signal_name> xor <signal_name>;
--    return <variable_name>; 
--  end <function_name>;

---- Example 2
--  function <function_name>  (signal <signal_name> : in <type_declaration>;
--                         signal <signal_name>   : in <type_declaration>  ) return <type_declaration> is
--  begin
--    if (<signal_name> = '1') then
--      return <signal_name>;
--    else
--      return 'Z';
--    end if;
--  end <function_name>;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;
 
end EthConstants;
