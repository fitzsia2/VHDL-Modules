---------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
---------------------------------------------------------------------------------
entity CRC_Ctrl is
   port(
      CLK_IN : in std_logic;
      COUNT_IN : in INTEGER;
      TXD : out std_logic_vector(3 downto 0) := (others => '0');
      LOADINIT_OUT : out std_logic := '0'; -- Initialize CRC generator
      START_CALC_OUT : out std_logic := '0'; -- Begin Calculating CRC
      DATA_VALID_OUT : out std_logic := '0'; -- Tell CRC generator the data is valid
      CLK_OUT: out std_logic := '0'; -- half the frequency of CLK_IN
      RCLK_OUT : out std_logic := '0'; -- Initiate read commands to memory
      DCLK_OUT : out std_logic := '0'; -- Send data to CRC generator
      DATA_IN : in std_logic_vector(63 downto 0) := X"0"; -- Accept data from memory
      RST_OUT : out std_logic := '0'); -- Restart CRC generator
end CRC_Ctrl;

---------------------------------------------------------------------------------
architecture Behavioral of CRC_Ctrl is


CONSTANT ETH_SFD1 : INTEGER := 11;
CONSTANT ETH_SFD2 : INTEGER := ETH_SFD1 + 1;
CONSTANT ETH_DESTADDR2 : INTEGER := ETH_SFD2 + 1;
CONSTANT ETH_DESTADDR1 : INTEGER := ETH_DESTADDR2 + 1;
CONSTANT ETH_DESTADDR4 : INTEGER := ETH_DESTADDR1 + 1;
CONSTANT ETH_DESTADDR3 : INTEGER := ETH_DESTADDR4 + 1;
CONSTANT ETH_DESTADDR6 : INTEGER := ETH_DESTADDR3 + 1;
CONSTANT ETH_DESTADDR5 : INTEGER := ETH_DESTADDR6 + 1;
CONSTANT ETH_DESTADDR8 : INTEGER := ETH_DESTADDR5 + 1;
CONSTANT ETH_DESTADDR7 : INTEGER := ETH_DESTADDR8 + 1;
CONSTANT ETH_DESTADDR10 : INTEGER := ETH_DESTADDR7 + 1;
CONSTANT ETH_DESTADDR9 : INTEGER := ETH_DESTADDR10 + 1;
CONSTANT ETH_DESTADDR12 : INTEGER := ETH_DESTADDR9 + 1;
CONSTANT ETH_DESTADDR11 : INTEGER := ETH_DESTADDR12 + 1;
CONSTANT ETH_SRCADDR2 : INTEGER := ETH_DESTADDR11 + 1;
CONSTANT ETH_SRCADDR1 : INTEGER := ETH_SRCADDR2 + 1;
CONSTANT ETH_SRCADDR4 : INTEGER := ETH_SRCADDR1 + 1;
CONSTANT ETH_SRCADDR3 : INTEGER := ETH_SRCADDR4 + 1;
CONSTANT ETH_SRCADDR6 : INTEGER := ETH_SRCADDR3 + 1;
CONSTANT ETH_SRCADDR5 : INTEGER := ETH_SRCADDR6 + 1;
CONSTANT ETH_SRCADDR8 : INTEGER := ETH_SRCADDR5 + 1;
CONSTANT ETH_SRCADDR7 : INTEGER := ETH_SRCADDR8 + 1;
CONSTANT ETH_SRCADDR10 : INTEGER := ETH_SRCADDR7 + 1;
CONSTANT ETH_SRCADDR9 : INTEGER := ETH_SRCADDR10 + 1;
CONSTANT ETH_SRCADDR12 : INTEGER := ETH_SRCADDR9 + 1;
CONSTANT ETH_SRCADDR11 : INTEGER := ETH_SRCADDR12 + 1;
CONSTANT ETH_TYPE2 : INTEGER := ETH_SRCADDR11 + 1;
CONSTANT ETH_TYPE1 : INTEGER := ETH_TYPE2 + 1;
CONSTANT ETH_TYPE4 : INTEGER := ETH_TYPE1 + 1;
CONSTANT ETH_TYPE3 : INTEGER := ETH_TYPE4 + 1;


   -- IPv4 Header Offsets

   -- 20Bytes
   -- 0  |0____.____|1____.____|2____.____|3____.____|
   -- 4  | Ver |Leng|Serv Type |     Total Length    |
   -- 8  |    Identification   |Flags|Fragment Offset|
   -- 12 |    TTL   | Protocol | Header Checksum     |
   -- 16 |             Source Address                |
   -- 20 |            Destination Address            |

   CONSTANT ETH_IPV4_IHL : INTEGER := ETH_TYPE3 + 1;
   CONSTANT ETH_IPV4_VER : INTEGER := ETH_IPV4_IHL + 1;
   CONSTANT ETH_IPV4_SRVTP2 : INTEGER := ETH_IPV4_VER + 1;
   CONSTANT ETH_IPV4_SRVTP1 : INTEGER := ETH_IPV4_SRVTP2 + 1;
   CONSTANT ETH_IPV4_LNG2 : INTEGER := ETH_IPV4_SRVTP1 + 1;
   CONSTANT ETH_IPV4_LNG1 : INTEGER := ETH_IPV4_LNG2 + 1;
   CONSTANT ETH_IPV4_LNG4 : INTEGER := ETH_IPV4_LNG1 + 1;
   CONSTANT ETH_IPV4_LNG3 : INTEGER := ETH_IPV4_LNG4 + 1;
   CONSTANT ETH_IPV4_ID2 : INTEGER := ETH_IPV4_LNG3 + 1;
   CONSTANT ETH_IPV4_ID1 : INTEGER := ETH_IPV4_ID2 + 1;
   CONSTANT ETH_IPV4_ID4 : INTEGER := ETH_IPV4_ID1 + 1;
   CONSTANT ETH_IPV4_ID3 : INTEGER := ETH_IPV4_ID4 + 1;
   CONSTANT ETH_IPV4_FRAGOFF1 : INTEGER := ETH_IPV4_ID3 + 1;
   CONSTANT ETH_IPV4_FLG : INTEGER := ETH_IPV4_FRAGOFF1 + 1;
   CONSTANT ETH_IPV4_FRAGOFF3 : INTEGER := ETH_IPV4_FLG + 1;
   CONSTANT ETH_IPV4_FRAGOFF2 : INTEGER := ETH_IPV4_FRAGOFF3 + 1;
   CONSTANT ETH_IPV4_LIVETIME2 : INTEGER := ETH_IPV4_FRAGOFF2 + 1;
   CONSTANT ETH_IPV4_LIVETIME1 : INTEGER := ETH_IPV4_LIVETIME2 + 1;
   CONSTANT ETH_IPV4_PROTOCOL2 : INTEGER := ETH_IPV4_LIVETIME1 + 1;
   CONSTANT ETH_IPV4_PROTOCOL1 : INTEGER := ETH_IPV4_PROTOCOL2 + 1;
   CONSTANT ETH_IPV4_HEADERCHKSM2 : INTEGER := ETH_IPV4_PROTOCOL1 + 1;
   CONSTANT ETH_IPV4_HEADERCHKSM1 : INTEGER := ETH_IPV4_HEADERCHKSM2 + 1;
   CONSTANT ETH_IPV4_HEADERCHKSM4 : INTEGER := ETH_IPV4_HEADERCHKSM1 + 1;
   CONSTANT ETH_IPV4_HEADERCHKSM3 : INTEGER := ETH_IPV4_HEADERCHKSM4 + 1;
   CONSTANT ETH_IPV4_SRCIP2 : INTEGER := ETH_IPV4_HEADERCHKSM3 + 1;
   CONSTANT ETH_IPV4_SRCIP1 : INTEGER := ETH_IPV4_SRCIP2 + 1;
   CONSTANT ETH_IPV4_SRCIP4 : INTEGER := ETH_IPV4_SRCIP1 + 1;
   CONSTANT ETH_IPV4_SRCIP3 : INTEGER := ETH_IPV4_SRCIP4 + 1;
   CONSTANT ETH_IPV4_SRCIP6 : INTEGER := ETH_IPV4_SRCIP3 + 1;
   CONSTANT ETH_IPV4_SRCIP5 : INTEGER := ETH_IPV4_SRCIP6 + 1;
   CONSTANT ETH_IPV4_SRCIP8 : INTEGER := ETH_IPV4_SRCIP5 + 1;
   CONSTANT ETH_IPV4_SRCIP7 : INTEGER := ETH_IPV4_SRCIP8 + 1;
   CONSTANT ETH_IPV4_DSTIP2 : INTEGER := ETH_IPV4_SRCIP7 + 1;
   CONSTANT ETH_IPV4_DSTIP1 : INTEGER := ETH_IPV4_DSTIP2 + 1;
   CONSTANT ETH_IPV4_DSTIP4 : INTEGER := ETH_IPV4_DSTIP1 + 1;
   CONSTANT ETH_IPV4_DSTIP3 : INTEGER := ETH_IPV4_DSTIP4 + 1;
   CONSTANT ETH_IPV4_DSTIP6 : INTEGER := ETH_IPV4_DSTIP3 + 1;
   CONSTANT ETH_IPV4_DSTIP5 : INTEGER := ETH_IPV4_DSTIP6 + 1;
   CONSTANT ETH_IPV4_DSTIP8 : INTEGER := ETH_IPV4_DSTIP5 + 1;
   CONSTANT ETH_IPV4_DSTIP7 : INTEGER := ETH_IPV4_DSTIP8 + 1;
   CONSTANT ETH_IPV4_PAYLOAD : INTEGER := ETH_IPV4_DSTIP7 + 1;


      -- UDP Header Offsets
      -- 8Bytes
      -- 0  |0____.____|1____.____|2____.____|3____.____|
      -- 4  |    Source Address   | Destination Address |
      -- 8  |        Length       |       Checksum      |
      CONSTANT ETH_IPV4_UDP_SRCADR2 : INTEGER := ETH_IPV4_DSTIP7 + 1;
      CONSTANT ETH_IPV4_UDP_SRCADR1 : INTEGER := ETH_IPV4_UDP_SRCADR2 + 1;
      CONSTANT ETH_IPV4_UDP_SRCADR4 : INTEGER := ETH_IPV4_UDP_SRCADR1 + 1;
      CONSTANT ETH_IPV4_UDP_SRCADR3 : INTEGER := ETH_IPV4_UDP_SRCADR4 + 1;
      CONSTANT ETH_IPV4_UDP_DSTADR2 : INTEGER := ETH_IPV4_UDP_SRCADR3 + 1;
      CONSTANT ETH_IPV4_UDP_DSTADR1 : INTEGER := ETH_IPV4_UDP_DSTADR2 + 1;
      CONSTANT ETH_IPV4_UDP_DSTADR4 : INTEGER := ETH_IPV4_UDP_DSTADR1 + 1;
      CONSTANT ETH_IPV4_UDP_DSTADR3 : INTEGER := ETH_IPV4_UDP_DSTADR4 + 1;
      CONSTANT ETH_IPV4_UDP_LENG2 : INTEGER   := ETH_IPV4_UDP_DSTADR3 + 1;
      CONSTANT ETH_IPV4_UDP_LENG1 : INTEGER   := ETH_IPV4_UDP_LENG2 + 1;
      CONSTANT ETH_IPV4_UDP_LENG4 : INTEGER   := ETH_IPV4_UDP_LENG1 + 1;
      CONSTANT ETH_IPV4_UDP_LENG3 : INTEGER   := ETH_IPV4_UDP_LENG4 + 1;
      CONSTANT ETH_IPV4_UDP_CHKSUM2 : INTEGER := ETH_IPV4_UDP_LENG3 + 1;
      CONSTANT ETH_IPV4_UDP_CHKSUM1 : INTEGER := ETH_IPV4_UDP_CHKSUM2 + 1;
      CONSTANT ETH_IPV4_UDP_CHKSUM4 : INTEGER := ETH_IPV4_UDP_CHKSUM1 + 1;
      CONSTANT ETH_IPV4_UDP_CHKSUM3 : INTEGER := ETH_IPV4_UDP_CHKSUM4 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N2 : INTEGER := ETH_IPV4_UDP_CHKSUM3 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N1 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N2 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N4 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N1  + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N3 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N4 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N6 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N3 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N5 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N6 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N8 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N5 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N7 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N8 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N10 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N7 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N9 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N10 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N12 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N9 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N11 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N12 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N14 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N11 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N13 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N14 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N16 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N13 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N15 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N16 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N18 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N15 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N17 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N18 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N20 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N17 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N19 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N20 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N22 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N19 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N21 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N22 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N24 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N21 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N23 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N24 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N26 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N23 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N25 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N26 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N28 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N25 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N27 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N28 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N30 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N27 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N29 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N30 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N32 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N29 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N31 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N32 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N34 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N31 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N33 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N34 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N36 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N33 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N35 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N36 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N38 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N35 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N37 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N38 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N40 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N37 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N39 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N40 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N42 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N39 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N41 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N42 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N44 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N41 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N43 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N44 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N46 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N43 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N45 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N46 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N48 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N45 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD_N47 : INTEGER := ETH_IPV4_UDP_PAYLOAD_N48 + 1;
      CONSTANT ETH_IPV4_UDP_PAYLOAD : INTEGER := ETH_IPV4_UDP_PAYLOAD_N47;
      
     
CONSTANT ETH_IPV4_DUP_ENDOFPAYLOAD : INTEGER := ETH_IPV4_UDP_PAYLOAD; -- = (ETH_IPV4_UDP_PAYLOAD) + (UDP Payload size)
CONSTANT ETH_IP_ENDOFPAYLOAD : INTEGER := ETH_IPV4_UDP_PAYLOAD; -- = (ETH_IPV4_UDP_PAYLOAD) + (UDP Payload size)
CONSTANT ETH_PAYLOAD : INTEGER := ETH_IPV4_UDP_PAYLOAD; -- Consider changing this to where CRC begins

CONSTANT ETH_CRC2 : INTEGER := ETH_IPV4_UDP_PAYLOAD + 1;
CONSTANT ETH_CRC1 : INTEGER := ETH_CRC2 + 1;
CONSTANT ETH_CRC4 : INTEGER := ETH_CRC1 + 1;
CONSTANT ETH_CRC3 : INTEGER := ETH_CRC4 + 1;
CONSTANT ETH_CRC6 : INTEGER := ETH_CRC3 + 1;
CONSTANT ETH_CRC5 : INTEGER := ETH_CRC6 + 1;
CONSTANT ETH_CRC8 : INTEGER := ETH_CRC5 + 1;
CONSTANT ETH_CRC7 : INTEGER := ETH_CRC8 + 1;

CONSTANT ETH_END_FRAME : INTEGER := ETH_CRC7 + 1;

CONSTANT ETH_FRAMEGAP : INTEGER := ETH_CRC7 + 24;

----------------------------------------
-- Ethernet frame constructors
----------------------------------------
-- Ethernet Header Constants
CONSTANT ETHPREAMBLE : STD_LOGIC_VECTOR := "1010";
CONSTANT SFD1 : STD_LOGIC_VECTOR := X"5";
CONSTANT SFD2 : STD_LOGIC_VECTOR := X"D";
CONSTANT BROADCAST : STD_LOGIC_VECTOR := X"F";
CONSTANT MAC_DESTADDR1 : STD_LOGIC_VECTOR := X"0";  -- 0 -- 00-1d-92-f3-31-53
CONSTANT MAC_DESTADDR2 : STD_LOGIC_VECTOR := X"0";  -- 0
CONSTANT MAC_DESTADDR3 : STD_LOGIC_VECTOR := X"1";  -- 1
CONSTANT MAC_DESTADDR4 : STD_LOGIC_VECTOR := X"D";  -- D
CONSTANT MAC_DESTADDR5 : STD_LOGIC_VECTOR := X"9";  -- 9
CONSTANT MAC_DESTADDR6 : STD_LOGIC_VECTOR := X"2";  -- 2
CONSTANT MAC_DESTADDR7 : STD_LOGIC_VECTOR := X"F";  -- F
CONSTANT MAC_DESTADDR8 : STD_LOGIC_VECTOR := X"3";  -- 3
CONSTANT MAC_DESTADDR9 : STD_LOGIC_VECTOR := X"3";  -- 3
CONSTANT MAC_DESTADDR10 : STD_LOGIC_VECTOR := X"1";  -- 1
CONSTANT MAC_DESTADDR11 : STD_LOGIC_VECTOR := X"5";  -- 5
CONSTANT MAC_DESTADDR12 : STD_LOGIC_VECTOR := X"3";  -- 3
CONSTANT MAC_SRCADDR1 : STD_LOGIC_VECTOR := X"A";  -- A -- A3-1C-6D-DF-B6-B6
CONSTANT MAC_SRCADDR2 : STD_LOGIC_VECTOR := X"3";  -- 3
CONSTANT MAC_SRCADDR3 : STD_LOGIC_VECTOR := X"1";  -- 1
CONSTANT MAC_SRCADDR4 : STD_LOGIC_VECTOR := X"C";  -- C
CONSTANT MAC_SRCADDR5 : STD_LOGIC_VECTOR := X"6";  -- 6
CONSTANT MAC_SRCADDR6 : STD_LOGIC_VECTOR := X"D";  -- D
CONSTANT MAC_SRCADDR7 : STD_LOGIC_VECTOR := X"D";  -- D
CONSTANT MAC_SRCADDR8 : STD_LOGIC_VECTOR := X"F";  -- F
CONSTANT MAC_SRCADDR9 : STD_LOGIC_VECTOR := X"B";  -- B
CONSTANT MAC_SRCADDR10 : STD_LOGIC_VECTOR := X"6"; -- 6
CONSTANT MAC_SRCADDR11 : STD_LOGIC_VECTOR := X"B"; -- B
CONSTANT MAC_SRCADDR12 : STD_LOGIC_VECTOR := X"6"; -- 6
CONSTANT ETHERTYPE1 : STD_LOGIC_VECTOR := X"0"; -- 0
CONSTANT ETHERTYPE2 : STD_LOGIC_VECTOR := X"8"; -- 8
CONSTANT ETHERTYPE3 : STD_LOGIC_VECTOR := X"0"; -- 0
CONSTANT ETHERTYPE4 : STD_LOGIC_VECTOR := X"0"; -- 0
CONSTANT CRC1 : STD_LOGIC_VECTOR := X"7"; -- bd890fc8 --> http://www.zorc.breitbandkatze.de/crc.html
CONSTANT CRC2 : STD_LOGIC_VECTOR := X"0"; -- d6fe9a4b --> Test bench
CONSTANT CRC3 : STD_LOGIC_VECTOR := X"7";
CONSTANT CRC4 : STD_LOGIC_VECTOR := X"0";
CONSTANT CRC5 : STD_LOGIC_VECTOR := X"A";
CONSTANT CRC6 : STD_LOGIC_VECTOR := X"D";
CONSTANT CRC7 : STD_LOGIC_VECTOR := X"F";
CONSTANT CRC8 : STD_LOGIC_VECTOR := X"C";

-- IPv4 Header Constants
CONSTANT IP_VER : STD_LOGIC_VECTOR := X"4";
CONSTANT IP_IHL : STD_LOGIC_VECTOR := X"5";
CONSTANT IP_SRVTP1 : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_SRVTP2 : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_LENG1 : STD_LOGIC_VECTOR := X"0"; -- = (20 Byte IP header) + (8 Byte UDP header) + (UDP payload) = 52
CONSTANT IP_LENG2 : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_LENG3 : STD_LOGIC_VECTOR := X"3";
CONSTANT IP_LENG4 : STD_LOGIC_VECTOR := X"4";
CONSTANT IP_ID : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_FLAGS : STD_LOGIC_VECTOR := X"4"; -- 11:7
CONSTANT IP_OFFSET : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_TTL1 : STD_LOGIC_VECTOR := X"F";
CONSTANT IP_TTL2 : STD_LOGIC_VECTOR := X"F";
CONSTANT IP_PROTOCOL1 : STD_LOGIC_VECTOR := X"1"; -- UDP Protocol ID
CONSTANT IP_PROTOCOL2 : STD_LOGIC_VECTOR := X"1";
CONSTANT IP_HDCHKSUM1 : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_HDCHKSUM2 : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_HDCHKSUM3 : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_HDCHKSUM4 : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_SRCIP1 : STD_LOGIC_VECTOR := X"C"; -- IP source is 192
CONSTANT IP_SRCIP2 : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_SRCIP3 : STD_LOGIC_VECTOR := X"A"; -- .168
CONSTANT IP_SRCIP4 : STD_LOGIC_VECTOR := X"8";
CONSTANT IP_SRCIP5 : STD_LOGIC_VECTOR := X"8"; -- .137
CONSTANT IP_SRCIP6 : STD_LOGIC_VECTOR := X"9";
CONSTANT IP_SRCIP7 : STD_LOGIC_VECTOR := X"7"; -- .120
CONSTANT IP_SRCIP8 : STD_LOGIC_VECTOR := X"8";
CONSTANT IP_DSTIP1 : STD_LOGIC_VECTOR := X"C"; -- IP destination is 192
CONSTANT IP_DSTIP2 : STD_LOGIC_VECTOR := X"0";
CONSTANT IP_DSTIP3 : STD_LOGIC_VECTOR := X"A"; -- .168
CONSTANT IP_DSTIP4 : STD_LOGIC_VECTOR := X"8";
CONSTANT IP_DSTIP5 : STD_LOGIC_VECTOR := X"8"; -- .137
CONSTANT IP_DSTIP6 : STD_LOGIC_VECTOR := X"9";
CONSTANT IP_DSTIP7 : STD_LOGIC_VECTOR := X"0"; -- .1
CONSTANT IP_DSTIP8 : STD_LOGIC_VECTOR := X"1";

-- UDP Header Constants
CONSTANT UDP_SRCADR1 : STD_LOGIC_VECTOR := X"0"; -- Least significant nibble
CONSTANT UDP_SRCADR2 : STD_LOGIC_VECTOR := X"A";
CONSTANT UDP_SRCADR3 : STD_LOGIC_VECTOR := X"0";
CONSTANT UDP_SRCADR4 : STD_LOGIC_VECTOR := X"A"; -- Most significant nibble
CONSTANT UDP_DSTADR1 : STD_LOGIC_VECTOR := X"0";
CONSTANT UDP_DSTADR2 : STD_LOGIC_VECTOR := X"C";
CONSTANT UDP_DSTADR3 : STD_LOGIC_VECTOR := X"0";
CONSTANT UDP_DSTADR4 : STD_LOGIC_VECTOR := X"0";
CONSTANT UDP_LENG1 : STD_LOGIC_VECTOR := X"0"; -- (8Byte header) + (24Byte payload) = 32
CONSTANT UDP_LENG2 : STD_LOGIC_VECTOR := X"0";
CONSTANT UDP_LENG3 : STD_LOGIC_VECTOR := X"2";
CONSTANT UDP_LENG4 : STD_LOGIC_VECTOR := X"0";
CONSTANT UDP_CHKSUM : STD_LOGIC_VECTOR := X"0"; -- 0
CONSTANT UDP_DATA_N1 : STD_LOGIC_VECTOR := X"1";
CONSTANT UDP_DATA_N2 : STD_LOGIC_VECTOR := X"2";
CONSTANT UDP_DATA_N3 : STD_LOGIC_VECTOR := X"3";
CONSTANT UDP_DATA_N4 : STD_LOGIC_VECTOR := X"4";
CONSTANT UDP_DATA_N5 : STD_LOGIC_VECTOR := X"5";
CONSTANT UDP_DATA_N6 : STD_LOGIC_VECTOR := X"6";
CONSTANT UDP_DATA_N7 : STD_LOGIC_VECTOR := X"7";
CONSTANT UDP_DATA_N8 : STD_LOGIC_VECTOR := X"8";
CONSTANT UDP_DATA_N9 : STD_LOGIC_VECTOR := X"9";
CONSTANT UDP_DATA_NA : STD_LOGIC_VECTOR := X"A";
CONSTANT UDP_DATA_NB : STD_LOGIC_VECTOR := X"B";
CONSTANT UDP_DATA_NC : STD_LOGIC_VECTOR := X"C";
CONSTANT UDP_DATA_ND : STD_LOGIC_VECTOR := X"D";
CONSTANT UDP_DATA_NE : STD_LOGIC_VECTOR := X"E";
CONSTANT UDP_DATA_NF : STD_LOGIC_VECTOR := X"F";
CONSTANT UDP_DATA_N0 : STD_LOGIC_VECTOR := X"0";

CONSTANT END_OF_TX1 : STD_LOGIC_VECTOR := "01101";
CONSTANT END_OF_TX2 : STD_LOGIC_VECTOR := "00111";

   signal Clk_DIV_16 : std_logic := '0';
   signal ClkOut_i : std_logic := '0';
   signal EthCounter_i : INTEGER := 0;
   
---------------------------------------------------------------------------------
-- Signal Assignments
--
begin
   CLK_OUT <= ClkOut_i;
   COUNT_OUT <= EthCounter_i;

---------------------------------------------------------------------------------
-- State Machine
--
--process( EthCounter_i )
--begin
--   if( EthCounter_i <= ETH_SFD1 ) then
--      TXD <= ETHPREAMBLE;
--   elsif( EthCounter_i < ETH_IPV4_UDP_PAYLOAD_N2 ) then -- N2 is the first byte
--      case EthCounter_i is
--      when ETH_SFD1 => TXD <= SFD1;
--      when ETH_SFD2 => TXD <= SFD2;
--      when ETH_DESTADDR1 => TXD <= MAC_DESTADDR1;
--      when ETH_DESTADDR2 => TXD <= MAC_DESTADDR2;
--      when ETH_DESTADDR3 => TXD <= MAC_DESTADDR3;
--      when ETH_DESTADDR4 => TXD <= MAC_DESTADDR4;
--      when ETH_DESTADDR5 => TXD <= MAC_DESTADDR5;
--      when ETH_DESTADDR6 => TXD <= MAC_DESTADDR6;
--      when ETH_DESTADDR7 => TXD <= MAC_DESTADDR7;
--      when ETH_DESTADDR8 => TXD <= MAC_DESTADDR8;
--      when ETH_DESTADDR9 => TXD <= MAC_DESTADDR9;
--      when ETH_DESTADDR10 => TXD <= MAC_DESTADDR10;
--      when ETH_DESTADDR11 => TXD <= MAC_DESTADDR11;
--      when ETH_DESTADDR12 => TXD <= MAC_DESTADDR12;
--      when ETH_SRCADDR1 => TXD <= MAC_SRCADDR1;
--      when ETH_SRCADDR2 => TXD <= MAC_SRCADDR2;
--      when ETH_SRCADDR3 => TXD <= MAC_SRCADDR3;
--      when ETH_SRCADDR4 => TXD <= MAC_SRCADDR4;
--      when ETH_SRCADDR5 => TXD <= MAC_SRCADDR5;
--      when ETH_SRCADDR6 => TXD <= MAC_SRCADDR6;
--      when ETH_SRCADDR7 => TXD <= MAC_SRCADDR7;
--      when ETH_SRCADDR8 => TXD <= MAC_SRCADDR8;
--      when ETH_SRCADDR9 => TXD <= MAC_SRCADDR9;
--      when ETH_SRCADDR10 => TXD <= MAC_SRCADDR10;
--      when ETH_SRCADDR11 => TXD <= MAC_SRCADDR11;
--      when ETH_SRCADDR12 => TXD <= MAC_SRCADDR12;
--      when ETH_TYPE1 => TXD <= ETHERTYPE1;
--      when ETH_TYPE2 => TXD <= ETHERTYPE2;
--      when ETH_TYPE3 => TXD <= ETHERTYPE3;
--      when ETH_TYPE4 => TXD <= ETHERTYPE4;
--      when ETH_IPV4_IHL => TXD <= IP_VER;
--      when ETH_IPV4_VER => TXD <= IP_IHL;
--      when ETH_IPV4_SRVTP1 => TXD <= IP_SRVTP1;
--      when ETH_IPV4_SRVTP2 => TXD <= IP_SRVTP2;
--      when ETH_IPV4_LNG1 => TXD <= IP_LENG1;
--      when ETH_IPV4_LNG2 => TXD <= IP_LENG2;
--      when ETH_IPV4_LNG3 => TXD <= IP_LENG3;
--      when ETH_IPV4_LNG4 => TXD <= IP_LENG4;
--      when ETH_IPV4_ID1 => TXD <= IP_ID;
--      when ETH_IPV4_ID2 => TXD <= IP_ID;
--      when ETH_IPV4_ID3 => TXD <= IP_ID;
--      when ETH_IPV4_ID4 => TXD <= IP_ID;
--      when ETH_IPV4_FLG => TXD <= IP_FLAGS;
--      when ETH_IPV4_FRAGOFF1 => TXD <= IP_OFFSET;
--      when ETH_IPV4_FRAGOFF2 => TXD <= IP_OFFSET;
--      when ETH_IPV4_FRAGOFF3 => TXD <= IP_OFFSET;
--      when ETH_IPV4_LIVETIME1 => TXD <= IP_TTL1;
--      when ETH_IPV4_LIVETIME2 => TXD <= IP_TTL2;
--      when ETH_IPV4_PROTOCOL1 => TXD <= IP_PROTOCOL1;
--      when ETH_IPV4_PROTOCOL2 => TXD <= IP_PROTOCOL2;
--      when ETH_IPV4_HEADERCHKSM1 => TXD <= IP_HDCHKSUM1;
--      when ETH_IPV4_HEADERCHKSM2 => TXD <= IP_HDCHKSUM2;
--      when ETH_IPV4_HEADERCHKSM3 => TXD <= IP_HDCHKSUM3;
--      when ETH_IPV4_HEADERCHKSM4 => TXD <= IP_HDCHKSUM4;
--      when ETH_IPV4_SRCIP1 => TXD <= IP_SRCIP1;
--      when ETH_IPV4_SRCIP2 => TXD <= IP_SRCIP2;
--      when ETH_IPV4_SRCIP3 => TXD <= IP_SRCIP3;
--      when ETH_IPV4_SRCIP4 => TXD <= IP_SRCIP4;
--      when ETH_IPV4_SRCIP5 => TXD <= IP_SRCIP5;
--      when ETH_IPV4_SRCIP6 => TXD <= IP_SRCIP6;
--      when ETH_IPV4_SRCIP7 => TXD <= IP_SRCIP7;
--      when ETH_IPV4_SRCIP8 => TXD <= IP_SRCIP8;
--      when ETH_IPV4_DSTIP1 => TXD <= IP_DSTIP1;
--      when ETH_IPV4_DSTIP2 => TXD <= IP_DSTIP2;
--      when ETH_IPV4_DSTIP3 => TXD <= IP_DSTIP3;
--      when ETH_IPV4_DSTIP4 => TXD <= IP_DSTIP4;
--      when ETH_IPV4_DSTIP5 => TXD <= IP_DSTIP5;
--      when ETH_IPV4_DSTIP6 => TXD <= IP_DSTIP6;
--      when ETH_IPV4_DSTIP7 => TXD <= IP_DSTIP7;
--      when ETH_IPV4_DSTIP8 => TXD <= IP_DSTIP8;
--      when ETH_IPV4_UDP_SRCADR1 => TXD <= UDP_SRCADR1;
--      when ETH_IPV4_UDP_SRCADR2 => TXD <= UDP_SRCADR2;
--      when ETH_IPV4_UDP_SRCADR3 => TXD <= UDP_SRCADR3;
--      when ETH_IPV4_UDP_SRCADR4 => TXD <= UDP_SRCADR4;
--      when ETH_IPV4_UDP_DSTADR1 => TXD <= UDP_DSTADR1;
--      when ETH_IPV4_UDP_DSTADR2 => TXD <= UDP_DSTADR2;
--      when ETH_IPV4_UDP_DSTADR3 => TXD <= UDP_DSTADR3;
--      when ETH_IPV4_UDP_DSTADR4 => TXD <= UDP_DSTADR4;
--      when ETH_IPV4_UDP_LENG1 => TXD <= UDP_LENG1;
--      when ETH_IPV4_UDP_LENG2 => TXD <= UDP_LENG2;
--      when ETH_IPV4_UDP_LENG3 => TXD <= UDP_LENG3;
--      when ETH_IPV4_UDP_LENG4 => TXD <= UDP_LENG4;
--      when ETH_IPV4_UDP_CHKSUM1 => TXD <= UDP_CHKSUM;
--      when ETH_IPV4_UDP_CHKSUM2 => TXD <= UDP_CHKSUM;
--      when ETH_IPV4_UDP_CHKSUM3 => TXD <= UDP_CHKSUM;
--      when ETH_IPV4_UDP_CHKSUM4 => TXD <= UDP_CHKSUM;
--      end case;
--   elsif( EthCounter_i > ETH_IPV4_UDP_CHKSUM3 and EthCounter_i <= ETH_IPV4_UDP_PAYLOAD ) then -- UDP Payload section
--      -- Load Camera Data Here
--   end if;
--end process;


---------------------------------------------------------------------------------
end Behavioral;

ARCHITECTURE txd_state of CRC_Ctrl is
begin
   with EthCounter_i select
      TXD <= "0000" when <= ETH_SFD1,
             "ZZZZ" when others;
end txd_state;


